module mux2(y,a,b,c);
input a;
input b;
input c;
output y;
assign y = (a&~c) | (b&c);
endmodule

module mux16to1(y,a,sel);
input [15:0] a;
input [3:0] sel;
wire [13:0] cables;
output y;

mux2 mux_1(cables[0],a[0],a[1],sel[0]);
mux2 mux_2(cables[1],a[2],a[3],sel[0]);
mux2 mux_3(cables[2],a[4],a[5],sel[0]);
mux2 mux_4(cables[3],a[6],a[7],sel[0]);
mux2 mux_5(cables[4],a[8],a[9],sel[0]);
mux2 mux_6(cables[5],a[10],a[11],sel[0]);
mux2 mux_7(cables[6],a[12],a[13],sel[0]);
mux2 mux_8(cables[7],a[14],a[15],sel[0]);

mux2 mux_9(cables[8],cables[0],cables[1],sel[1]);
mux2 mux_10(cables[9],cables[2],cables[3],sel[1]);
mux2 mux_11(cables[10],cables[4],cables[5],sel[1]);
mux2 mux_12(cables[11],cables[6],cables[7],sel[1]);

mux2 mux_13(cables[12],cables[8],cables[9],sel[2]);
mux2 mux_14(cables[13],cables[10],cables[11],sel[2]);

mux2 mux_15(y,cables[12],cables[13],sel[3]);

endmodule

module mux16to1_tb;
reg [15:0] a;
reg [3:0] sel;
wire y;
mux16to1 prueba(y,a,sel);
initial begin
a[0]=1;a[1]=0;a[2]=0; a[3] = 0; a[4] = 0; a[5] = 0; a[6] = 0; a[7] = 0; a[8] = 0; a[9] = 0; a[10] = 0; a[11] = 0; a[12] = 0; a[13] = 0; a[14] = 0; a[15] = 0; sel[3] = 0; sel[2] = 0;sel[1] = 0; sel[0] = 0;
#1
a[0]=0;a[1]=1;a[2]=0; a[3] = 0; a[4] = 0; a[5] = 0; a[6] = 0; a[7] = 0; a[8] = 0; a[9] = 0; a[10] = 0; a[11] = 0; a[12] = 0; a[13] = 0; a[14] = 0; a[15] = 0; sel[3] = 0; sel[2] = 0;sel[1] = 0; sel[0] = 1;
#1
a[0]=0;a[1]=0;a[2]=1; a[3] = 0; a[4] = 0; a[5] = 0; a[6] = 0; a[7] = 0; a[8] = 0; a[9] = 0; a[10] = 0; a[11] = 0; a[12] = 0; a[13] = 0; a[14] = 0; a[15] = 0; sel[3] = 0; sel[2] = 0;sel[1] = 1; sel[0] = 0;
#1
a[0]=0;a[1]=0;a[2]=0; a[3] = 1; a[4] = 0; a[5] = 0; a[6] = 0; a[7] = 0; a[8] = 0; a[9] = 0; a[10] = 0; a[11] = 0; a[12] = 0; a[13] = 0; a[14] = 0; a[15] = 0; sel[3] = 0; sel[2] = 0;sel[1] = 1; sel[0] = 1;
#1
a[0]=0;a[1]=0;a[2]=0; a[3] = 0; a[4] = 1; a[5] = 0; a[6] = 0; a[7] = 0; a[8] = 0; a[9] = 0; a[10] = 0; a[11] = 0; a[12] = 0; a[13] = 0; a[14] = 0; a[15] = 0; sel[3] = 0; sel[2] = 1;sel[1] = 0; sel[0] = 0;
#1
a[0]=0;a[1]=0;a[2]=0; a[3] = 0; a[4] = 0; a[5] = 1; a[6] = 0; a[7] = 0; a[8] = 0; a[9] = 0; a[10] = 0; a[11] = 0; a[12] = 0; a[13] = 0; a[14] = 0; a[15] = 0; sel[3] = 0; sel[2] = 1;sel[1] = 0; sel[0] = 1;
#1
a[0]=0;a[1]=0;a[2]=0; a[3] = 0; a[4] = 0; a[5] = 0; a[6] = 1; a[7] = 0; a[8] = 0; a[9] = 0; a[10] = 0; a[11] = 0; a[12] = 0; a[13] = 0; a[14] = 0; a[15] = 0; sel[3] = 0; sel[2] = 1;sel[1] = 1; sel[0] = 0;
#1
a[0]=0;a[1]=0;a[2]=0; a[3] = 0; a[4] = 0; a[5] = 0; a[6] = 0; a[7] = 1; a[8] = 0; a[9] = 0; a[10] = 0; a[11] = 0; a[12] = 0; a[13] = 0; a[14] = 0; a[15] = 0; sel[3] = 0; sel[2] = 1;sel[1] = 1; sel[0] = 1;
#1
a[0]=0;a[1]=0;a[2]=0; a[3] = 0; a[4] = 0; a[5] = 0; a[6] = 0; a[7] = 0; a[8] = 1; a[9] = 0; a[10] = 0; a[11] = 0; a[12] = 0; a[13] = 0; a[14] = 0; a[15] = 0; sel[3] = 1; sel[2] = 0;sel[1] = 0; sel[0] = 0;
#1
a[0]=0;a[1]=0;a[2]=0; a[3] = 0; a[4] = 0; a[5] = 0; a[6] = 0; a[7] = 0; a[8] = 0; a[9] = 1; a[10] = 0; a[11] = 0; a[12] = 0; a[13] = 0; a[14] = 0; a[15] = 0; sel[3] = 1; sel[2] = 0;sel[1] = 0; sel[0] = 1;
#1
a[0]=0;a[1]=0;a[2]=0; a[3] = 0; a[4] = 0; a[5] = 0; a[6] = 0; a[7] = 0; a[8] = 0; a[9] = 0; a[10] = 1; a[11] = 0; a[12] = 0; a[13] = 0; a[14] = 0; a[15] = 0; sel[3] = 1; sel[2] = 0;sel[1] = 1; sel[0] = 0;
#1
a[0]=0;a[1]=0;a[2]=0; a[3] = 0; a[4] = 0; a[5] = 0; a[6] = 0; a[7] = 0; a[8] = 0; a[9] = 0; a[10] = 0; a[11] = 1; a[12] = 0; a[13] = 0; a[14] = 0; a[15] = 0; sel[3] = 1; sel[2] = 0;sel[1] = 1; sel[0] = 1;
#1
a[0]=0;a[1]=0;a[2]=0; a[3] = 0; a[4] = 0; a[5] = 0; a[6] = 0; a[7] = 0; a[8] = 0; a[9] = 0; a[10] = 0; a[11] = 0; a[12] = 1; a[13] = 0; a[14] = 0; a[15] = 0; sel[3] = 1; sel[2] = 1;sel[1] = 0; sel[0] = 0;
#1
a[0]=0;a[1]=0;a[2]=0; a[3] = 0; a[4] = 0; a[5] = 0; a[6] = 0; a[7] = 0; a[8] = 0; a[9] = 0; a[10] = 0; a[11] = 0; a[12] = 0; a[13] = 1; a[14] = 0; a[15] = 0; sel[3] = 1; sel[2] = 1;sel[1] = 0; sel[0] = 1;
#1
a[0]=0;a[1]=0;a[2]=0; a[3] = 0; a[4] = 0; a[5] = 0; a[6] = 0; a[7] = 0; a[8] = 0; a[9] = 0; a[10] = 0; a[11] = 0; a[12] = 0; a[13] = 0; a[14] = 1; a[15] = 0; sel[3] = 1; sel[2] = 1;sel[1] = 1; sel[0] = 0;
#1
a[0]=0;a[1]=0;a[2]=0; a[3] = 0; a[4] = 0; a[5] = 0; a[6] = 0; a[7] = 0; a[8] = 0; a[9] = 0; a[10] = 0; a[11] = 0; a[12] = 0; a[13] = 0; a[14] = 0; a[15] = 1; sel[3] = 1; sel[2] = 1;sel[1] = 1; sel[0] = 1;
#1
    $finish;
end
initial begin
    $monitor("%2d\t a0 = %b\t a1 = %b\t a2 = %b\ta3 = %b\ta4 = %b\ta5 = %b\ta6 = %b\ta7 = %b\ta8 = %b\ta9 = %b\ta10 = %b\ta11 = %b\ta12 = %b\ta13 = %b\ta14 = %b\ta15 = %b\ty = %b\t",$time,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],y);
end
endmodule
