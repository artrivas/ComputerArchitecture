module tristate(y,a,enable);
input a;
input enable;
output y;

endmodule
