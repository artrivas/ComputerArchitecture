module behavioral_srlatch(Q,Qn,S,R);
input S,R;
output Q,Qn;

endmodule
